--entity validate is
--	generic
--	(
--		<name>	: <type>  :=	<default_value>;
--		...
--		<name>	: <type>  :=	<default_value>
--	);
--
--
--	port
--	(
--		-- Input ports
--		<name>	: in  <type>;
--		<name>	: in  <type> := <default_value>;
--
--		-- Inout ports
--		<name>	: inout <type>;
--
--		-- Output ports
--		<name>	: out <type>;
--		<name>	: out <type> := <default_value>
--	);
--end validate;
