library ieee;
use ieee.std_logic_1164.all;

entity reg is
  generic (
    N : integer := 4
  );
  port (
    clk : in std_logic;
    data_in : in std_logic_vector(N-1 downto 0);
    data_out : out std_logic_vector(N-1 downto 0);
    load : in std_logic; -- Write enable
    clear : in std_logic
  );
end reg;

architecture rtl of reg is

begin
  -- Your code here!
  process (Clk, load, clear) 
  variable temp : std_logic_vector(N-1 downto 0);
  begin 
	if (clear = '1') 	then
		temp := "0000";
	elsif Clk'EVENT AND Clk = '1' and load = '1' then
		temp := data_in;
	end if;
	data_out <= temp;
	
  end process;
end rtl;
